module main

import ss 

fn main() {
	mut app := ss.new_app();
	app.run()!;
}
